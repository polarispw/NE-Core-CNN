module conv1_buf #(parameter WIDTH = 28, HEIGHT = 28, DATA_BITS = 8)(
   input clk,
   input rst_n,
   input [DATA_BITS - 1:0] data_in,
   output reg [DATA_BITS - 1:0] data_out_0, data_out_1, data_out_2, data_out_3, data_out_4,
   data_out_5, data_out_6, data_out_7, data_out_8, data_out_9,
   data_out_10, data_out_11, data_out_12, data_out_13, data_out_14,
   data_out_15, data_out_16, data_out_17, data_out_18, data_out_19,
   data_out_20, data_out_21, data_out_22, data_out_23, data_out_24,
   output reg valid_out_buf
 );

 localparam FILTER_SIZE = 5;

 reg [DATA_BITS - 1:0] buffer [0:WIDTH * FILTER_SIZE - 1];
 reg [DATA_BITS - 1:0] buf_idx;
 reg [4:0] w_idx, h_idx;
 reg [2:0] buf_flag;  // 0 ~ 4
 reg state;

 always @(posedge clk) begin
   if(~rst_n) begin
     buf_idx <= -1;
     w_idx <= 0;
     h_idx <= 0;
     buf_flag <= 0;
     state <= 0;
     valid_out_buf <= 0;
     data_out_0 <= 12'bx;
     data_out_1 <= 12'bx;
     data_out_2 <= 12'bx;
     data_out_3 <= 12'bx;
     data_out_4 <= 12'bx;
     data_out_5 <= 12'bx;
     data_out_6 <= 12'bx;
     data_out_7 <= 12'bx;
     data_out_8 <= 12'bx;
     data_out_9 <= 12'bx;
     data_out_10 <= 12'bx;
     data_out_11 <= 12'bx;
     data_out_12 <= 12'bx;
     data_out_13 <= 12'bx;
     data_out_14 <= 12'bx;
     data_out_15 <= 12'bx;
     data_out_16 <= 12'bx;
     data_out_17 <= 12'bx;
     data_out_18 <= 12'bx;
     data_out_19 <= 12'bx;
     data_out_20 <= 12'bx;
     data_out_21 <= 12'bx;
     data_out_22 <= 12'bx;
     data_out_23 <= 12'bx;
     data_out_24 <= 12'bx;
   end 
   //创建一个28×5的buffer，当加载完140个数据后，从第一排开始继续更新数据
   
   else begin
      buf_idx <= buf_idx + 1;
      if(buf_idx == WIDTH * FILTER_SIZE - 1) begin // buffer size = 140 = 28(w) * 5(h)
        buf_idx <= 0;
      end
      
      buffer[buf_idx] <= data_in;  // data input
      
      // Wait until first 140 input data filled in buffer
      if(!state) begin                               //state为0时进行数据加载，为1时进行卷积操作
        if(buf_idx == WIDTH * FILTER_SIZE - 1) begin
          state <= 1'b1;                            //加载完140个数据后，state变1，开始进行以下卷积操作
        end
      end 

      else begin // valid state
        w_idx <= w_idx + 1'b1; // move right

        if(w_idx == WIDTH - FILTER_SIZE + 1) begin
          valid_out_buf <= 1'b0; // unvalid area    //第一排卷积操作结束，让valid_out_buf变0，从而使后面的max池化层停止操作；等待这一排的后几个数据更新完毕再变回1
        end 
        
        else if(w_idx == WIDTH - 1) begin        
          buf_flag <= buf_flag + 1'b1;              //第一排数据更新完毕后，更改buf_flag模式，此时的buffer第一排相当于实际28×28数据的第6排；以此类推
          if(buf_flag == FILTER_SIZE - 1) begin
            buf_flag <= 0;                          //当28×5的5行全部更新完毕，相当于又重新回到最开始加载完140个数据的模式，buf_flag变回最开始的模式
          end
          w_idx <= 0;                                //5行更新完毕后，5×28的buffer的行索引w_idx重新归0

          if(h_idx == HEIGHT - FILTER_SIZE) begin  // done 1 input read -> 28 * 28
            h_idx <= 0;                            //28×28整个输入数据的行索引，在所有卷积操作完成后归0
            state <= 1'b0;							//在所有卷积操作完毕后state归0，停止卷积操作
          end 
          
          h_idx <= h_idx + 1'b1;
        end 

        else if(w_idx == 0) begin
          valid_out_buf <= 1'b1; // start valid area    //每卷积并更新完一行数据后valid_out_buf变1传递到max池化层，开始池化操作
        end

        // Buffer Selection -> 5 * 5
        if(buf_flag == 3'd0) begin
          data_out_0 <= buffer[w_idx];
          data_out_1 <= buffer[w_idx + 1];
          data_out_2 <= buffer[w_idx + 2];
          data_out_3 <= buffer[w_idx + 3];
          data_out_4 <= buffer[w_idx + 4];

          data_out_5 <= buffer[w_idx + WIDTH];
          data_out_6 <= buffer[w_idx + 1 + WIDTH];
          data_out_7 <= buffer[w_idx + 2 + WIDTH];
          data_out_8 <= buffer[w_idx + 3 + WIDTH];
          data_out_9 <= buffer[w_idx + 4 + WIDTH];

          data_out_10 <= buffer[w_idx + WIDTH * 2];
          data_out_11 <= buffer[w_idx + 1 + WIDTH * 2];
          data_out_12 <= buffer[w_idx + 2 + WIDTH * 2];
          data_out_13 <= buffer[w_idx + 3 + WIDTH * 2];
          data_out_14 <= buffer[w_idx + 4 + WIDTH * 2];

          data_out_15 <= buffer[w_idx + WIDTH * 3];
          data_out_16 <= buffer[w_idx + 1 + WIDTH * 3];
          data_out_17 <= buffer[w_idx + 2 + WIDTH * 3];
          data_out_18 <= buffer[w_idx + 3 + WIDTH * 3];
          data_out_19 <= buffer[w_idx + 4 + WIDTH * 3];

          data_out_20 <= buffer[w_idx + WIDTH * 4];
          data_out_21 <= buffer[w_idx + 1 + WIDTH * 4];
          data_out_22 <= buffer[w_idx + 2 + WIDTH * 4];
          data_out_23 <= buffer[w_idx + 3 + WIDTH * 4];
          data_out_24 <= buffer[w_idx + 4 + WIDTH * 4];
        end else if(buf_flag == 3'd1) begin
          data_out_0 <= buffer[w_idx + WIDTH];
          data_out_1 <= buffer[w_idx + 1 + WIDTH];
          data_out_2 <= buffer[w_idx + 2 + WIDTH];
          data_out_3 <= buffer[w_idx + 3 + WIDTH];
          data_out_4 <= buffer[w_idx + 4 + WIDTH];

          data_out_5 <= buffer[w_idx + WIDTH * 2];
          data_out_6 <= buffer[w_idx + 1 + WIDTH * 2];
          data_out_7 <= buffer[w_idx + 2 + WIDTH * 2];
          data_out_8 <= buffer[w_idx + 3 + WIDTH * 2];
          data_out_9 <= buffer[w_idx + 4 + WIDTH * 2];

          data_out_10 <= buffer[w_idx + WIDTH * 3];
          data_out_11 <= buffer[w_idx + 1 + WIDTH * 3];
          data_out_12 <= buffer[w_idx + 2 + WIDTH * 3];
          data_out_13 <= buffer[w_idx + 3 + WIDTH * 3];
          data_out_14 <= buffer[w_idx + 4 + WIDTH * 3];

          data_out_15 <= buffer[w_idx + WIDTH * 4];
          data_out_16 <= buffer[w_idx + 1 + WIDTH * 4];
          data_out_17 <= buffer[w_idx + 2 + WIDTH * 4];
          data_out_18 <= buffer[w_idx + 3 + WIDTH * 4];
          data_out_19 <= buffer[w_idx + 4 + WIDTH * 4];

          data_out_20 <= buffer[w_idx];
          data_out_21 <= buffer[w_idx + 1];
          data_out_22 <= buffer[w_idx + 2];
          data_out_23 <= buffer[w_idx + 3];
          data_out_24 <= buffer[w_idx + 4];
        end else if(buf_flag == 3'd2) begin
          data_out_0 <= buffer[w_idx + WIDTH * 2];
          data_out_1 <= buffer[w_idx + 1 + WIDTH * 2];
          data_out_2 <= buffer[w_idx + 2 + WIDTH * 2];
          data_out_3 <= buffer[w_idx + 3 + WIDTH * 2];
          data_out_4 <= buffer[w_idx + 4 + WIDTH * 2];

          data_out_5 <= buffer[w_idx + WIDTH * 3];
          data_out_6 <= buffer[w_idx + 1 + WIDTH * 3];
          data_out_7 <= buffer[w_idx + 2 + WIDTH * 3];
          data_out_8 <= buffer[w_idx + 3 + WIDTH * 3];
          data_out_9 <= buffer[w_idx + 4 + WIDTH * 3];

          data_out_10 <= buffer[w_idx + WIDTH * 4];
          data_out_11 <= buffer[w_idx + 1 + WIDTH * 4];
          data_out_12 <= buffer[w_idx + 2 + WIDTH * 4];
          data_out_13 <= buffer[w_idx + 3 + WIDTH * 4];
          data_out_14 <= buffer[w_idx + 4 + WIDTH * 4];

          data_out_15 <= buffer[w_idx];
          data_out_16 <= buffer[w_idx + 1];
          data_out_17 <= buffer[w_idx + 2];
          data_out_18 <= buffer[w_idx + 3];
          data_out_19 <= buffer[w_idx + 4];

          data_out_20 <= buffer[w_idx + WIDTH];
          data_out_21 <= buffer[w_idx + 1 + WIDTH];
          data_out_22 <= buffer[w_idx + 2 + WIDTH];
          data_out_23 <= buffer[w_idx + 3 + WIDTH];
          data_out_24 <= buffer[w_idx + 4 + WIDTH];
        end else if(buf_flag == 3'd3) begin
          data_out_0 <= buffer[w_idx + WIDTH * 3];
          data_out_1 <= buffer[w_idx + 1 + WIDTH * 3];
          data_out_2 <= buffer[w_idx + 2 + WIDTH * 3];
          data_out_3 <= buffer[w_idx + 3 + WIDTH * 3];
          data_out_4 <= buffer[w_idx + 4 + WIDTH * 3];

          data_out_5 <= buffer[w_idx + WIDTH * 4];
          data_out_6 <= buffer[w_idx + 1 + WIDTH * 4];
          data_out_7 <= buffer[w_idx + 2 + WIDTH * 4];
          data_out_8 <= buffer[w_idx + 3 + WIDTH * 4];
          data_out_9 <= buffer[w_idx + 4 + WIDTH * 4];

          data_out_10 <= buffer[w_idx];
          data_out_11 <= buffer[w_idx + 1];
          data_out_12 <= buffer[w_idx + 2];
          data_out_13 <= buffer[w_idx + 3];
          data_out_14 <= buffer[w_idx + 4];

          data_out_15 <= buffer[w_idx + WIDTH];
          data_out_16 <= buffer[w_idx + 1 + WIDTH];
          data_out_17 <= buffer[w_idx + 2 + WIDTH];
          data_out_18 <= buffer[w_idx + 3 + WIDTH];
          data_out_19 <= buffer[w_idx + 4 + WIDTH];

          data_out_20 <= buffer[w_idx + WIDTH * 2];
          data_out_21 <= buffer[w_idx + 1 + WIDTH * 2];
          data_out_22 <= buffer[w_idx + 2 + WIDTH * 2];
          data_out_23 <= buffer[w_idx + 3 + WIDTH * 2];
          data_out_24 <= buffer[w_idx + 4 + WIDTH * 2];      
        end else if(buf_flag == 3'd4) begin
          data_out_0 <= buffer[w_idx + WIDTH * 4];
          data_out_1 <= buffer[w_idx + 1 + WIDTH * 4];
          data_out_2 <= buffer[w_idx + 2 + WIDTH * 4];
          data_out_3 <= buffer[w_idx + 3 + WIDTH * 4];
          data_out_4 <= buffer[w_idx + 4 + WIDTH * 4];

          data_out_5 <= buffer[w_idx];
          data_out_6 <= buffer[w_idx + 1];
          data_out_7 <= buffer[w_idx + 2];
          data_out_8 <= buffer[w_idx + 3];
          data_out_9 <= buffer[w_idx + 4];

          data_out_10 <= buffer[w_idx + WIDTH];
          data_out_11 <= buffer[w_idx + 1 + WIDTH];
          data_out_12 <= buffer[w_idx + 2 + WIDTH];
          data_out_13 <= buffer[w_idx + 3 + WIDTH];
          data_out_14 <= buffer[w_idx + 4 + WIDTH];

          data_out_15 <= buffer[w_idx + WIDTH * 2];
          data_out_16 <= buffer[w_idx + 1 + WIDTH * 2];
          data_out_17 <= buffer[w_idx + 2 + WIDTH * 2];
          data_out_18 <= buffer[w_idx + 3 + WIDTH * 2];
          data_out_19 <= buffer[w_idx + 4 + WIDTH * 2];

          data_out_20 <= buffer[w_idx + WIDTH * 3];
          data_out_21 <= buffer[w_idx + 1 + WIDTH * 3];
          data_out_22 <= buffer[w_idx + 2 + WIDTH * 3];
          data_out_23 <= buffer[w_idx + 3 + WIDTH * 3];
          data_out_24 <= buffer[w_idx + 4 + WIDTH * 3];   
        end
      end
   end
 end
endmodule

